`timescale 1ns / 1ps

//AXI ST VIP�ӿڵĶ�Ŀ����

module ikun_multi_target_detect #(
    parameter   IMG_HDISP   =   1280,   //ͼ��ˮƽ�ֱ���
    parameter   IMG_VDISP   =   720 ,   //ͼ����ֱ�ֱ���
    parameter   MIN_DIST    =   30      //��Ŀ������뾶
)
(
    input                       clk,
    input                       rst_n,
        
    input   wire                s_axis_video_tdata,
    input   wire                s_axis_video_tvalid,
    output  reg                 s_axis_video_tready,
    input   wire                s_axis_video_tlast,
    input   wire                s_axis_video_tuser,

	output	reg	    [44:0]		target_pos_out [15:0],	// {Flag,ymax[43:33],xmax[32:22],ymin[21:11],xmin[10:0]}
    output  reg     [ 3:0]      target_num_out,         //����Ŀ����Ŀ      
    output  reg                 target_pos_valid        //Ŀ��ϲ���ɣ����Ŀ���ַ��Ч
    );
    
reg         video_in_data   ;
reg         video_in_valid  ; 
reg         video_in_ready  ;
reg         video_in_last   ;
reg         video_in_user   ;

reg         video_data_dly  ;
reg         video_valid_dly ; 
reg         video_last_dly  ;
reg         video_user_dly  ;

//////////////////////////////////////////////////////////step 1
//register axis input, insert bubble cycles

always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        s_axis_video_tready <=  1'b0;
        
        video_in_data       <=  1'b0;
        video_in_valid      <=  1'b0;
        video_in_last       <=  1'b0;
        video_in_user       <=  1'b0;
    end
    else begin
        if(s_axis_video_tready) begin
            s_axis_video_tready <=  !s_axis_video_tvalid;
            
            video_in_data       <=  s_axis_video_tdata;
            video_in_valid      <=  s_axis_video_tvalid;
            video_in_last       <=  s_axis_video_tlast;
            video_in_user       <=  s_axis_video_tuser;
        end
        else if(video_in_ready) begin
            s_axis_video_tready <=  1'b1;
            
            video_in_valid      <=  1'b0;
        end
    end
end

//////////////////////////////////////////////////////////step 2
//delay for a clock cycle

always @(posedge clk or negedge rst_n) begin
    if(!rst_n) begin       
        video_data_dly      <=  1'b0;
        video_valid_dly     <=  1'b0;
        video_last_dly      <=  1'b0;
        video_user_dly      <=  1'b0;
    end
    else begin
        video_data_dly      <=  video_in_valid && video_in_ready && video_in_data;
        video_valid_dly     <=  video_in_valid && video_in_ready                 ;
        video_last_dly      <=  video_in_valid && video_in_ready && video_in_last;
        video_user_dly      <=  video_in_valid && video_in_ready && video_in_user;
    end
end


//------------------------------------------
//��������ͷ����ͼ�����������
reg [10:0] video_in_x_cnt;    
reg [10:0] video_in_y_cnt;    

always @ (posedge clk or negedge rst_n) begin
    if(!rst_n) begin
        video_in_x_cnt <= 11'd0;
        video_in_y_cnt <= 11'd0;
    end
    else if(video_in_valid && video_in_ready) begin
        if(video_in_last) begin
            video_in_x_cnt <= 11'd0;   
            video_in_y_cnt <= video_in_y_cnt + 1'b1;   
        end
        else if(video_in_user) begin
            video_in_x_cnt <= 11'd0;       
            video_in_y_cnt <= 11'd0;
        end
        else begin
            video_in_x_cnt <= video_in_x_cnt + 1'b1;       
        end
    end  
end

//------------------------------------------
//�Ĵ�����
reg [10:0]  x_cnt_r;
reg [10:0]  y_cnt_r;

always@(posedge clk or negedge rst_n) begin
	if(!rst_n)  begin
        x_cnt_r <= 11'd0;
		y_cnt_r <= 11'd0;
	end
	else begin
		x_cnt_r <= video_in_x_cnt;
        y_cnt_r <= video_in_y_cnt;
	end
end

//------------------------------------------
// {Flag,ymax[43:33],xmax[32:22],ymin[21:11],xmin[10:0]}
reg  [44:0]	target_pos		        [15:0] ;	//�Ĵ�����˶�Ŀ��ı߽� 

wire [15:0] target_flag;				        //��Ŀ�����Ч��־					 
wire [10:0] target_boarder_left 	[15:0] ;	//��Ŀ�����/��/��/�±߽�  
wire [10:0] target_boarder_right 	[15:0] ;								 
wire [10:0] target_boarder_top		[15:0] ;								 
wire [10:0] target_boarder_bottom	[15:0] ;	

wire [10:0] target_left 	        [15:0] ;	//��Ŀ������ķ�Χ  
wire [10:0] target_right 	        [15:0] ;								 
wire [10:0] target_top		        [15:0] ;								 
wire [10:0] target_bottom	        [15:0] ;	

generate
genvar i; 
	for(i=0; i<16; i = i+1) begin: list
		assign target_flag[i]           =  target_pos[i][44]; 

		assign target_boarder_bottom[i] =  target_pos[i][43:33];	//�±߽����������
		assign target_boarder_right[i]  =  target_pos[i][32:22];	//�ұ߽����������
		assign target_boarder_top[i]    =  target_pos[i][21:11];	//�ϱ߽����������
		assign target_boarder_left[i]   =  target_pos[i][10: 0];	//��߽����������
        
		assign target_bottom[i] =  (target_pos[i][43:33] < IMG_VDISP-1 - MIN_DIST  ) ? (target_pos[i][43:33] + MIN_DIST) : IMG_VDISP-1;	//�±߽����������
		assign target_right[i]  =  (target_pos[i][32:22] < IMG_HDISP-1 - MIN_DIST  ) ? (target_pos[i][32:22] + MIN_DIST) : IMG_HDISP-1;	//�ұ߽����������
		assign target_top[i]    =  (target_pos[i][21:11] > 11'd0       + MIN_DIST  ) ? (target_pos[i][21:11] - MIN_DIST) : 11'd0;		//�ϱ߽����������
		assign target_left[i]   =  (target_pos[i][10: 0] > 11'd0       + MIN_DIST  ) ? (target_pos[i][10: 0] - MIN_DIST) : 11'd0;		//��߽����������

	end
endgenerate

//------------------------------------------
//��Ⲣ���Ŀ����Ҫ��������ʱ�� 
integer j ;
reg [ 3:0] target_cnt;
reg [15:0] new_target_flag;		//��⵽��Ŀ���ͶƱ��	 

always@(posedge clk or negedge rst_n) begin
	if(!rst_n) begin
		//��ʼ�����˶�Ŀ��ı߽�Ϊ0
		for(j=0; j<16; j = j+1) begin	
			target_pos[j] <= {1'b0,11'd0,11'd0,11'd0,11'd0};
		end
		new_target_flag	<= 16'd0;
		target_cnt 		<= 4'd0;
	end
		//��һ֡��ʼ���г�ʼ��
	else if(video_in_valid && video_in_ready && video_in_user)begin  
		for(j=0; j<16; j = j+1) begin	
			target_pos[j] <= {1'b0,11'd0,11'd0,11'd0,11'd0};
		end
		new_target_flag	<= 16'd0;
		target_cnt 		<= 4'd0;
	end  
	else begin 
	//------------------------------------------
    //��һ��ʱ�����ڣ��ҳ����Ϊ�˶�Ŀ������ص㣬���˶�Ŀ���б��е�Ԫ�ؽ���ͶƱ���ж��Ƿ�Ϊȫ�µ��˶�Ŀ��
		if(video_in_valid && video_in_ready && video_in_data) begin		 
			for(j=0; j<16; j = j+1) begin
				if(target_flag[j] == 1'b0) begin		//�˶�Ŀ���б��е�������Ч�����Ԫ��ͶƱ�϶�����ĻҶ�Ϊ�µ����ֵ					
					new_target_flag[j] <= 1'b1; 
				end	
				else begin								//�˶�Ŀ���б��е�������Ч�����жϵ�ǰ�����Ƿ����ڸ�Ԫ��������
					if((video_in_x_cnt < target_left[j]) || (video_in_x_cnt > target_right[j])
                            ||(video_in_y_cnt < target_top[j])||(video_in_y_cnt > target_bottom[j])) begin 
						new_target_flag[j] <= 1'b1;		//���������볬��Ŀ������Χ��ͶƱ�϶�Ϊ�µ�Ŀ��
					end	
					else begin
						new_target_flag[j] <= 1'b0;		//�����϶�Ϊ�µ�Ŀ��	
					end
				end
			end
		end
		else begin
            new_target_flag	<= 16'd0;					//�������ص㲻���˶�Ŀ�� 
        end  
		
        //------------------------------------------
		//�ڶ���ʱ�����ڣ�����ͶƱ���������ѡ���ݸ��µ��˶�Ŀ���б���
		if(video_valid_dly && video_data_dly) begin 
			if(new_target_flag == 16'hffff)begin  		//ȫƱͨ������־�ų����µ��˶�Ŀ�� 
				target_pos[target_cnt] <= {1'b1,y_cnt_r,x_cnt_r,y_cnt_r,x_cnt_r};
				target_cnt <= target_cnt + 1'b1;
			end	
			else if (new_target_flag > 16'd0)begin		//���ֱ����Ϊ�˶�Ŀ������ص㣬���������˶�Ŀ���б���ĳ��Ԫ�ص�������
			
				for(j=0; j<16; j = j+1) begin	       	//�����˶�Ŀ���б���չ���и�Ԫ�ص�����Χ
				
					if(new_target_flag[j] == 1'b0) begin //δͶƱ�϶�Ϊ��Ŀ���Ԫ�أ���ʾ��ǰ����λ������������
					
						target_pos[j][44] 		<= 1'b1; 
						
						if(x_cnt_r < target_pos[j][10: 0] )		//��X����С����߽磬����X������չΪ��߽�
							target_pos[j][10: 0] <= x_cnt_r ;
							
						if(x_cnt_r > target_pos[j][32:22] )		//��X��������ұ߽磬����X������չΪ�ұ߽�
							target_pos[j][32:22] <=	x_cnt_r ;
							
						if(y_cnt_r < target_pos[j][21:11] )		//��Y����С���ϱ߽磬����Y������չΪ�ϱ߽�
							target_pos[j][21:11] <=	y_cnt_r ;
							
						if(y_cnt_r > target_pos[j][43:33] )		//��Y��������±߽磬����Y������չΪ�±߽�
							target_pos[j][43:33] <=	y_cnt_r ;

					end
				end
				
			end  
		end
	end 
end 

/////////////////////////////////////////
//һ֡ͳ�ƽ����󣬼Ĵ�������
integer k;

reg [ 3:0] repet_target_cnt;    //�����ų��ظ���Ŀ��
reg [ 3:0] check_target_cnt;    //�����ų��ظ���Ŀ��
reg [ 3:0] valid_target_cnt;    //������Ч��Ŀ����
reg [ 3:0] delete_repet_state;  //״̬�������ڲ��Ҳ�ɾ���ظ�Ŀ��

reg	[44:0] target_pos_reg[15:0];//��ʱ�Ĵ������

always@(posedge clk or negedge rst_n)
begin
	if(!rst_n) begin
		for(k=0; k<16; k = k+1) begin	
			target_pos_out[k] <=  {1'b0,11'd0,11'd0,11'd0,11'd0};
			target_pos_reg[k] <=  {1'b0,11'd0,11'd0,11'd0,11'd0};
		end
        
        repet_target_cnt    <= 4'd0;
        check_target_cnt    <= 4'd0;
        valid_target_cnt    <= 4'd0;
        target_pos_valid    <= 1'b0;
        delete_repet_state  <= 4'd0;
        
        target_num_out      <= 4'd0;
        video_in_ready      <= 1'b1;
	end
	else begin
        case(delete_repet_state)
            4'd0: begin
                if((x_cnt_r == IMG_HDISP - 1) && (y_cnt_r == IMG_VDISP - 1))begin   //һ֡ͳ�ƽ���������Ĵ������㣬��ʼ���Ҳ�ɾ���ظ�Ŀ��
                    for(k=0; k<16; k = k+1) begin	
                        target_pos_out[k] <= {1'b0,11'd0,11'd0,11'd0,11'd0};
                        target_pos_reg[k] <= target_pos[k]; //�Ĵ��Ŀ����
                    end
                    
                    repet_target_cnt    <= 4'd0;            //�ӵ�0��Ŀ�꿪ʼ�ų�
                    check_target_cnt    <= 4'd1;            //�ɵ�1Ŀ�꿪ʼ�Ƚϣ�0Ŀ�겻�غ��Լ��Ƚϣ�
                    valid_target_cnt    <= 4'd0;
                    target_pos_valid    <= 1'b0;
                    delete_repet_state  <= 4'd1;
                    
                    video_in_ready      <= 1'b0;
                end
            end
    
            4'd1: begin
                if(target_pos_reg[repet_target_cnt][44] == 1'b0) begin    //�����ǰĿ���FLAG��־λΪ0��������Ŀ��������    
                    target_pos_valid    <= 1'b1;
                    delete_repet_state  <= 4'd0;
                    
                    target_num_out      <= valid_target_cnt; //�Ĵ����պϲ�֮���Ŀ����Ŀ
                    video_in_ready      <= 1'b1;
                end
                else if(target_pos_reg[check_target_cnt][44] == 1'b0) begin    //����Ƚ�Ŀ���FLAG��־λΪ0����ǰĿ�������    
                    delete_repet_state  <= 4'd2;
                end
                else begin  //Ŀ����Ч�����������Ŀ��Ƚϣ��ж��Ƿ����ص�����
                
                    //û���ص�����������һĿ������Ƚ�
                    if((target_pos_reg[repet_target_cnt][10: 0] > target_pos_reg[check_target_cnt][32:22]) ||       //��߽�����ұ߽�
                        (target_pos_reg[repet_target_cnt][32:22] < target_pos_reg[check_target_cnt][10: 0]) ||      //�ұ߽�С����߽�
                            (target_pos_reg[repet_target_cnt][21:11] > target_pos_reg[check_target_cnt][43:33]) ||  //�ϱ߽�����±߽�
                                (target_pos_reg[repet_target_cnt][43:33] < target_pos_reg[check_target_cnt][21:11]) //�±߽�С���ϱ߽�
                                    ) begin   
                        if(check_target_cnt < 4'd15) begin  //�����Ƚ���һ��Ŀ��
                            check_target_cnt    <= check_target_cnt + 1'b1;
                            delete_repet_state  <= 4'd1;
                        end
                        else begin
                            delete_repet_state  <= 4'd2;    //�Ƚϵ����һ��Ŀ�꣬��ǰĿ�������
                        end    
                    end
                    //���ص����򣬽���ǰĿ�������ϲ����Ƚ�Ŀ���У�ͬʱ�ų�����ǰĿ��
                    else begin                           
						if( target_pos_reg[repet_target_cnt][10: 0] <  target_pos_reg[check_target_cnt][10: 0] )		//��X����С����߽磬����X������չΪ��߽�
                            target_pos_reg[check_target_cnt][10: 0] <= target_pos_reg[repet_target_cnt][10: 0] ;
							
						if( target_pos_reg[repet_target_cnt][32:22] >  target_pos_reg[check_target_cnt][32:22] )		//��X��������ұ߽磬����X������չΪ�ұ߽�
							target_pos_reg[check_target_cnt][32:22] <= target_pos_reg[repet_target_cnt][32:22] ;
							
						if( target_pos_reg[repet_target_cnt][21:11]  < target_pos_reg[check_target_cnt][21:11] )		//��Y����С���ϱ߽磬����Y������չΪ�ϱ߽�
							target_pos_reg[check_target_cnt][21:11] <= target_pos_reg[repet_target_cnt][21:11]  ;
							
						if( target_pos_reg[repet_target_cnt][43:33] >  target_pos_reg[check_target_cnt][43:33] )		//��Y��������±߽磬����Y������չΪ�±߽�
							target_pos_reg[check_target_cnt][43:33] <= target_pos_reg[repet_target_cnt][43:33] ;

                        if(repet_target_cnt < 4'd14) begin      //�����ų���һ��Ŀ��
                            repet_target_cnt    <= repet_target_cnt + 1'b1;
                            check_target_cnt    <= repet_target_cnt + 4'd2;
                            delete_repet_state  <= 4'd1;
                        end
                        else begin
                            repet_target_cnt    <= repet_target_cnt + 1'b1; //���һ��Ŀ��ֱ����� 
                            delete_repet_state  <= 4'd2;
                        end
                    end
                end
            end
          
            4'd2: begin //Ŀ������ɣ�û���ظ�Ŀ�꣬����Ŀ��д�����յ�����ӿ�
                target_pos_out[valid_target_cnt] <= target_pos_reg[repet_target_cnt];
                
                valid_target_cnt        <= valid_target_cnt + 1'b1; 
                
                if(repet_target_cnt < 4'd14) begin //�����һ��Ŀ��
                    repet_target_cnt    <= repet_target_cnt + 1'b1; //���ֵΪ14
                    check_target_cnt    <= repet_target_cnt + 4'd2; //���ֵΪ15
                    delete_repet_state  <= 4'd1;    //�����ų�
                end
                else if(repet_target_cnt == 4'd14) begin   //��һ��Ŀ��Ϊ���һ��Ŀ�꣬���ü�飬ֱ�����
                    repet_target_cnt    <= repet_target_cnt + 1'b1; //���һ��Ŀ��Ϊ15
                    delete_repet_state  <= 4'd2;    //ֱ�����
                end
                else begin
                    target_pos_valid    <= 1'b1;    //����Ŀ��Ƚ����
                    delete_repet_state  <= 4'd0;
                    
                    target_num_out      <= valid_target_cnt; //�Ĵ����պϲ�֮���Ŀ����Ŀ
                    
                    video_in_ready      <= 1'b1;
                end
            end
    
        endcase
        
    end
end
    
endmodule
